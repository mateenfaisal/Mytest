module added (a, b, c)
input a,b;
output c;
endmodule
